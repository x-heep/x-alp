package core_v_mcu_pkg;



endpackage : core_v_mcu_pkg
