module cpu_subsystem (
    input logic clk_i,
    input logic rst_ni
);
    
    cva6 #(
        
    ) cpu_inst (

    );

endmodule
