package x_alp_pkg;

endpackage : x_alp_pkg
